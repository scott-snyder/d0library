 UPGRADED D0   BIPOLAR PULSE   DET C=4.7NF
 0.6268
 0.1200
 0.000D+00  0.000D+00 .             X             .             .             .
 1.000D-07  0.000D+00 .             *+            .             .             .
 2.000D-07  1.196D-04 .             *     +       .             .             .
 3.000D-07  1.730D-02 .             . *          +.             .             .
 4.000D-07  6.069D-02 .             .       *     .   +         .             .
 5.000D-07  1.005D-01 .             .             *       +     .             .
 6.000D-07  1.197D-01 .             .             .  *      +   .             .
 7.000D-07  1.139D-01 .             .             . *        +  .             .
 8.000D-07  8.402D-02 .             .           * .           + .             .
 9.000D-07  4.371D-02 .             .     *       .          +  .             .
 1.000D-06  4.641D-03 .             .*            .          +  .             .
 1.100D-06 -2.744D-02 .         *   .             .          +  .             .
 1.200D-06 -4.916D-02 .      *      .             .          +  .             .
 1.300D-06 -6.060D-02 .     *       .             .          +  .             .
 1.400D-06 -6.396D-02 .    *        .             .          +  .             .
 1.500D-06 -6.150D-02 .    *        .             .          +  .             .
 1.600D-06 -5.554D-02 .     *       .             .          +  .             .
 1.700D-06 -4.798D-02 .      *      .             .          +  .             .
 1.800D-06 -4.006D-02 .       *     .             .          +  .             .
 1.900D-06 -3.258D-02 .        *    .             .          +  .             .
 2.000D-06 -2.598D-02 .         *   .             .          +  .             .
 2.100D-06 -2.038D-02 .          *  .             .          +  .             .
 2.200D-06 -1.579D-02 .           * .             .          +  .             .
 2.300D-06 -1.211D-02 .           * .             .          +  .             .
 2.400D-06 -9.210D-03 .            *.             .          +  .             .
 2.500D-06 -6.955D-03 .            *.             .          +  .             .
 2.600D-06 -5.219D-03 .            *.             .          +  .             .
 2.700D-06 -3.894D-03 .            *.             .          +  .             .
 2.800D-06 -2.892D-03 .             *             .          +  .             .
 2.900D-06 -2.139D-03 .             *             .          +  .             .
 3.000D-06 -1.574D-03 .             *             .          +  .             .
 3.100D-06 -1.154D-03 .             *             .          +  .             .
 3.200D-06 -8.420D-04 .             *             .          +  .             .
 3.400D-06 -4.459D-04 .             *             .         +   .             .
 3.600D-06 -2.338D-04 .             *             .         +   .             .
 3.800D-06 -1.213D-04 .             *             .         +   .             .
 4.000D-06 -5.897D-05 .             *             .         +   .             .
 4.200D-06 -2.441D-05 .             *             .         +   .             .
 4.400D-06 -1.825D-05 .             *             .         +   .             .
 4.600D-06 -7.831D-06 .             *             .         +   .             .
 4.800D-06  1.094D-06 .             *             .         +   .             .
 5.000D-06  3.941D-06 .             *             .         +   .             .
 5.200D-06  4.082D-06 .             *             .         +   .             .
 5.400D-06  6.226D-06 .             *             .         +   .             .
 5.600D-06  7.588D-06 .             *             .         +   .             .
 5.800D-06 -2.819D-07 .             *             .         +   .             .
 6.000D-06  6.833D-07 .             *             .         +   .             .
 6.200D-06  5.733D-06 .             *             .         +   .             .
 6.400D-06  3.192D-07 .             *             .         +   .             .
