 D0 ORIGINAL ELECTRONICS     CDET=4.7 NF$                            
 2.200
 0.750
 0.000D+00  0.000D+00 *             +             .             .             .
 2.000D-07  3.154D-05 *             .+            .             .             .
 4.000D-07  3.040D-02 . *           .    +        .             .             .
 6.000D-07  1.220D-01 .        *    .         +   .             .             .
 8.000D-07  2.461D-01 .             .  *          .+            .             .
 1.000D-06  3.698D-01 .             .           * .   +         .             .
 1.200D-06  4.781D-01 .             .             .    *+       .             .
 1.400D-06  5.662D-01 .             .             .      +    * .             .
 1.600D-06  6.345D-01 .             .             .       +     . *           .
 1.800D-06  6.857D-01 .             .             .        +    .     *       .
 2.000D-06  7.229D-01 .             .             .         +   .        *    .
 2.200D-06  7.490D-01 .             .             .         +   .         *   .
 2.400D-06  7.668D-01 .             .             .         +   .           * .
 2.600D-06  7.781D-01 .             .             .         +   .           * .
 3.000D-06  7.879D-01 .             .             .         +   .            *.
 4.000D-06  7.770D-01 .             .             .         +   .           * .
 6.000D-06  7.232D-01 .             .             .         +   .        *    .
 8.000D-06  6.689D-01 .             .             .         *   .+            .
 1.000D-05  6.174D-01 .             .             . *  +        .             .
 2.000D-05  4.040D-01 .             .X            .             .             .
 3.000D-05  2.492D-01 .             .             +      *      .             .
 4.000D-05  1.378D-01 .             .    * +      .             .             .
 5.000D-05  5.862D-02 .       *    +.             .             .             .
 5.400D-05  3.411D-02 .    *    +   .             .             .             .
 5.800D-05  1.276D-02 . *     +     .             .             .             .
 6.000D-05  3.232D-03 *     +       .             .             .             .
 6.200D-05 -5.680D-03 .             .           * .    +        .             .
 6.400D-05 -1.384D-02 .             .         *   .   +         .             .
 6.600D-05 -2.143D-02 .             .       *     .  +          .             .
 6.800D-05 -2.843D-02 .             .     *       .+            .             .
 7.000D-05 -3.487D-02 .             .   *         .+            .             .
 7.500D-05 -4.887D-02 .             *        +    .             .             .
 8.000D-05 -6.032D-02 .          *  .  +          .             .             .
 9.000D-05 -7.655D-02 .      X      .             .             .             .
 1.000D-04 -8.614D-02 .   *        +.             .             .             .
 1.100D-04 -9.090D-02 .  *    +     .             .             .             .
 1.200D-04 -9.241D-02 . * +         .             .             .             .
 1.300D-04 -9.154D-02 .     *       .             +             .             .
 1.400D-04 -8.910D-02 .       *     .          +  .             .             .
 1.500D-04 -8.566D-02 .         *   .       +     .             .             .
 1.600D-04 -8.153D-02 .            *.    +        .             .             .
 1.700D-04 -7.704D-02 .             . X           .             .             .
 1.800D-04 -7.242D-02 .            +.    *        .             .             .
 1.900D-04 -6.776D-02 .          +  .        *    .             .             .
 2.000D-04 -6.326D-02 .        +    .           * .             .             .
 2.100D-04 -5.881D-02 .      +      .             .*            .             .
 2.200D-04 -5.462D-02 .    +        .             .   *         .             .
 2.300D-04 -5.063D-02 .   +         .             .      *      .             .
 2.400D-04 -4.686D-02 . +           .             .        *    .             .
