  UPGRADED D0  FAST UNIPOLAR PULSE  DET C=1NF
  0.6300 
  0.318
  8.000E-08     0.000E+00   3.554E-03
  1.200E-07     0.000E+00   4.356E-02
  2.000E-07     4.717E-08   1.745E-01
  2.400E-07     8.224E-04   2.541E-01
  2.600E-07     3.163E-03   2.874E-01
  2.800E-07     8.048E-03   3.181E-01
  3.000E-07     1.609E-02   3.473E-01
  3.200E-07     2.755E-02   3.749E-01
  3.400E-07     4.262E-02   4.016E-01
  3.600E-07     6.136E-02   4.330E-01
  3.800E-07     8.356E-02   4.700E-01
  4.000E-07     1.085E-01   5.112E-01
  4.200E-07     1.353E-01   5.529E-01
  4.400E-07     1.629E-01   5.946E-01
  4.600E-07     1.905E-01   6.379E-01
  4.800E-07     2.170E-01   6.822E-01
  5.000E-07     2.417E-01   7.249E-01
  5.200E-07     2.636E-01   7.624E-01
  5.400E-07     2.821E-01   7.945E-01
  5.600E-07     2.969E-01   8.227E-01
  5.800E-07     3.078E-01   8.481E-01
  6.000E-07     3.149E-01   8.698E-01
  6.200E-07     3.180E-01   8.860E-01
  6.400E-07     3.174E-01   8.983E-01
  6.600E-07     3.134E-01   9.086E-01
  6.800E-07     3.062E-01   9.187E-01
  7.000E-07     2.961E-01   9.274E-01
  7.200E-07     2.835E-01   9.338E-01
  7.400E-07     2.686E-01   9.384E-01
  7.600E-07     2.518E-01   9.423E-01
  7.800E-07     2.336E-01   9.463E-01
  8.000E-07     2.143E-01   9.486E-01
  8.200E-07     1.943E-01   9.489E-01
  8.400E-07     1.740E-01   9.475E-01
  8.800E-07     1.341E-01   9.440E-01
  9.200E-07     9.712E-02   9.379E-01
  1.000E-06     3.917E-02   9.259E-01
  1.080E-06     5.491E-03   9.202E-01
  1.160E-06    -8.820E-03   9.186E-01
  1.240E-06    -1.142E-02   9.180E-01
  1.320E-06    -8.478E-03   9.179E-01
  1.400E-06    -4.199E-03   9.186E-01
  1.480E-06    -9.561E-04   9.192E-01
  1.560E-06     6.091E-04   9.191E-01
  1.640E-06     9.373E-04   9.188E-01
  1.720E-06     6.649E-04   9.185E-01
  1.800E-06     2.086E-04   9.183E-01
  1.880E-06    -2.043E-04   9.180E-01
  2.000E-06    -1.0000-04   9.175E-01
