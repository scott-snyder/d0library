 UPGRADED D0   UNIPOLAR PULSE   DET C=4.7NF
 1.0220
 0.3568
 0.000D+00  0.000D+00 .             X             .             .             .
 1.000D-07  0.000D+00 .             X             .             .             .
 2.000D-07  8.303D-09 .             * +           .             .             .
 3.000D-07  1.421D-03 .             *    +        .             .             .
 4.000D-07  1.551D-02 .             .*       +    .             .             .
 5.000D-07  5.561D-02 .             .   *         +             .             .
 6.000D-07  1.226D-01 .             .        *    .    +        .             .
 7.000D-07  2.037D-01 .             .             *        +    .             .
 8.000D-07  2.799D-01 .             .             .     *    +  .             .
 9.000D-07  3.341D-01 .             .             .        *  + .             .
 1.000D-06  3.568D-01 .             .             .          *+ .             .
 1.100D-06  3.479D-01 .             .             .         * + .             .
 1.200D-06  3.137D-01 .             .             .       *   + .             .
 1.300D-06  2.635D-01 .             .             .   *       + .             .
 1.400D-06  2.070D-01 .             .             *          +  .             .
 1.500D-06  1.523D-01 .             .          *  .          +  .             .
 1.600D-06  1.045D-01 .             .      *      .          +  .             .
 1.700D-06  6.640D-02 .             .    *        .          +  .             .
 1.800D-06  3.829D-02 .             .  *          .          +  .             .
 1.900D-06  1.920D-02 .             .*            .          +  .             .
 2.000D-06  7.387D-03 .             .*            .          +  .             .
 2.100D-06  9.096D-04 .             *             .          +  .             .
 2.200D-06 -2.011D-03 .             *             .          +  .             .
 2.300D-06 -2.808D-03 .             *             .          +  .             .
 2.400D-06 -2.519D-03 .             *             .          +  .             .
 2.500D-06 -1.821D-03 .             *             .          +  .             .
 2.600D-06 -1.101D-03 .             *             .          +  .             .
 2.700D-06 -5.430D-04 .             *             .          +  .             .
 2.800D-06 -1.993D-04 .             *             .          +  .             .
 2.900D-06 -5.262D-05 .             *             .          +  .             .
 3.000D-06 -5.494D-05 .             *             .          +  .             .
 3.100D-06 -1.525D-04 .             *             .          +  .             .
 3.200D-06 -2.983D-04 .             *             .          +  .             .
 3.400D-06 -6.076D-04 .             *             .          +  .             .
 3.600D-06 -8.386D-04 .             *             .          +  .             .
 3.800D-06 -9.685D-04 .             *             .          +  .             .
 4.000D-06 -1.027D-03 .             *             .          +  .             .
 4.200D-06 -1.045D-03 .             *             .          +  .             .
 4.400D-06 -1.044D-03 .             *             .          +  .             .
 4.600D-06 -1.044D-03 .             *             .          +  .             .
 4.800D-06 -1.041D-03 .             *             .          +  .             .
 5.000D-06 -1.035D-03 .             *             .          +  .             .
 5.200D-06 -1.035D-03 .             *             .          +  .             .
 5.400D-06 -1.043D-03 .             *             .          +  .             .
 5.600D-06 -1.051D-03 .             *             .          +  .             .
 5.800D-06 -1.050D-03 .             *             .          +  .             .
 6.000D-06 -1.041D-03 .             *             .          +  .             .
 6.200D-06 -1.037D-03 .             *             .          +  .             .
 6.400D-06 -1.040D-03 .             *             .          +  .             .
